----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:43:03 07/21/2015 
-- Design Name: 
-- Module Name:    fsmc_glue - A_fsmc_glue 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.std_logic_misc.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity fsmc2bram_sync is
  Generic (
    AW_FSMC : positive;     -- total FSMC address width
    DW : positive;          -- data witdth
    AW_SLAVE : positive     -- actually used address lines starts from
  );
	Port (
    clk : in std_logic; -- extenal clock generated by FSMC bus
    mmu_int : out std_logic;
    
    A : in STD_LOGIC_VECTOR (AW_FSMC-1 downto 0);
    D : inout STD_LOGIC_VECTOR (DW-1 downto 0);
    NWE : in STD_LOGIC;
    NOE : in STD_LOGIC;
    NCE : in STD_LOGIC;
    
    bram_a   : out STD_LOGIC_VECTOR (AW_SLAVE-1 downto 0);
    bram_di  : in  STD_LOGIC_VECTOR (DW-1 downto 0);
    bram_do  : out STD_LOGIC_VECTOR (DW-1 downto 0);
    bram_ce  : out STD_LOGIC;
    bram_we  : out STD_LOGIC_VECTOR (0 downto 0);
    bram_clk : out std_logic
  );
  
end fsmc2bram_sync;



-----------------------------------------------------------------------------

architecture beh of fsmc2bram_sync is

  type state_t is (IDLE, ADSET, RECEIVE, TRANSMIT);
  signal state : state_t := IDLE;
  signal a_cnt : std_logic_vector(AW_SLAVE-1 downto 0) := (others => '0');
  signal data_reg_fsmc2bram : std_logic_vector(DW-1 downto 0) := (others => '0');
  signal data_reg_bram2fsmc : std_logic_vector(DW-1 downto 0) := (others => '0'); 
  
begin

  -- connect permanent signals
  bram_clk <= clk;
  bram_a   <= a_cnt;
  
  -- coonect 3-state data bus
  --D <= bram_di when (NCE = '0' and NOE = '0') else (others => 'Z');
  --bram_do <= D;
  D <= data_reg_bram2fsmc when (NCE = '0' and NOE = '0') else (others => 'Z');
  bram_do <= data_reg_fsmc2bram;
  bram_we <= "1" when (state = RECEIVE) else "0";
  bram_ce <= '1' when (state = RECEIVE or state = TRANSMIT) else '0';
  
  --
  --
  --
  mmu_process : process(clk) is
  begin
    if rising_edge(clk) then
      if (NCE = '0') then
        mmu_int <= or_reduce(A(AW_FSMC-1 downto AW_SLAVE));
      else
        mmu_int <= '0';
      end if;
    end if;
  end process;
  
  --
  --
  --
  fsmc_state_process : process(clk) is
    variable latcnt : std_logic_vector(1 downto 0) := (others => '0');
    variable tx_cycle : boolean := false;
  begin
    if rising_edge(clk) then
      if NCE = '1' then
        state <= IDLE;
        latcnt := (others => '0');
      else
        case state is
        when IDLE =>
          a_cnt <= A(AW_SLAVE-1 downto 0);
          if (NWE = '0') then
            latcnt := "10";
            tx_cycle := false;
          else
            latcnt := "11";
            tx_cycle := true;
          end if;
          state <= ADSET;

        when ADSET =>
          latcnt := latcnt - 1;
          if (latcnt = "000") then
            if tx_cycle then
              state <= TRANSMIT;
            else
              state <= RECEIVE;
            end if;
          end if;
          
        when TRANSMIT =>
          a_cnt <= a_cnt + 1;
          data_reg_bram2fsmc <= bram_di;
          
        when RECEIVE =>
          a_cnt <= a_cnt + 1;
          data_reg_fsmc2bram <= D;

        end case;
      end if; -- NCE
    end if; -- clk
  end process;


 
end beh;




